-- Insert Control Circuit (probably a FSM) Here