-- Insert top-level entity here